library verilog;
use verilog.vl_types.all;
entity shuma_vlg_vec_tst is
end shuma_vlg_vec_tst;
