library verilog;
use verilog.vl_types.all;
entity speed_ctrl_vlg_vec_tst is
end speed_ctrl_vlg_vec_tst;
