library verilog;
use verilog.vl_types.all;
entity lev_ctl_vlg_vec_tst is
end lev_ctl_vlg_vec_tst;
