module music_mem (
  input   wire            clk,
  input   wire            rst_n,
  
  input   wire    [9:0]   cnt,   // 10位输入
  
  output  reg     [4:0]   music
);

  // 1024×5位 ROM (32×1024位 = 4KB)
  reg [4:0] note_rom [0:1023];
  
  // 音符定义（根据lev_ctl.v的编码）
  parameter SIL = 5'd0;   // 静音
  //低音
  parameter LOW_C  = 5'd1;   // 01_001 = 低音Do
  parameter LOW_D  = 5'd2;   // 01_010 = 低音Re
  parameter LOW_E  = 5'd3;   // 01_011 = 低音Mi
  parameter LOW_F  = 5'd4;   // 01_100 = 低音Fa
  parameter LOW_G  = 5'd5;   // 01_101 = 低音Sol 
  parameter LOW_A  = 5'd6;   // 01_110 = 低音La  
  parameter LOW_B  = 5'd7;   // 01_111 = 低音Si
  // 中音
  parameter MID_C = 5'd9;   // 中音Do (10_001)
  parameter MID_D = 5'd10;  // 中音Re (10_010)
  parameter MID_E = 5'd11;  // 中音Mi (10_011)
  parameter MID_F = 5'd12;  // 中音Fa (10_100)
  parameter MID_G = 5'd13;  // 中音Sol (101_101)
  parameter MID_A = 5'd14;  // 中音La (10_110)
  parameter MID_B = 5'd15;  // 中音Si (10_111)
  // 高音
  parameter HIGH_C = 5'd17; // 高音Do (11_001)
  parameter HIGH_D = 5'd18; // 高音Re (11_010)
  parameter HIGH_E = 5'd19; // 高音Mi (11_011)
  parameter HIGH_F = 5'd20; // 高音Fa (11_100)
  parameter HIGH_G = 5'd21; // 高音Sol(11_101)
  parameter HIGH_A = 5'd22; // 高音La (11_110)
  parameter HIGH_B = 5'd23; // 高音Si (11_111)
  
  
  parameter HIGH_C2 = 5'd25; // 超高音Do
  
  // 初始化ROM
  integer i; 
  
  initial begin
    // 初始化为静音（0）
    for (i = 0; i < 1024; i = i + 1) begin
      note_rom[i] = SIL;
    end
   
//歌唱祖国	
    // ====== 第一首歌(地址 0-511) ======
    note_rom[0]    = LOW_G;
    note_rom[1]    = LOW_G;
    note_rom[2]    = LOW_G;
    note_rom[3]    = LOW_G;
    note_rom[4]    = MID_C;
    note_rom[5]    = MID_C;
    note_rom[6]    = MID_C;
    note_rom[7]    = MID_C;
    note_rom[8]    = LOW_G;
    note_rom[9]    = LOW_G;
    note_rom[10]   = LOW_G;
    note_rom[11]   = LOW_G;
    note_rom[12]   = MID_E;
    note_rom[13]   = MID_E;
    note_rom[14]   = MID_E;
    note_rom[15]   = MID_E;
    note_rom[16]   = MID_C;
    note_rom[17]   = MID_C;
    note_rom[18]   = MID_C;
    note_rom[19]   = MID_C;
    note_rom[20]   = MID_G;
    note_rom[21]   = MID_G;
    note_rom[22]   = MID_G;
    note_rom[23]   = MID_G;
    note_rom[24]   = MID_G;
    note_rom[25]   = MID_A;
    note_rom[26]   = MID_A;
    note_rom[27]   = MID_A;
    note_rom[28]   = MID_G;
    note_rom[29]   = MID_G;
    note_rom[30]   = MID_G;
    note_rom[31]   = MID_G;
    note_rom[32]   = SIL;
    note_rom[33]   = MID_G;
    note_rom[34]   = MID_G;
    note_rom[35]   = MID_G;
    note_rom[36]   = MID_G;
    note_rom[37]   = MID_G;
    note_rom[38]   = MID_G;
    note_rom[39]   = HIGH_C;
    note_rom[40]   = HIGH_C;
    note_rom[41]   = HIGH_C;
    note_rom[42]   = HIGH_C;
    note_rom[43]   = HIGH_C;
    note_rom[44]   = HIGH_C;
    note_rom[45]   = HIGH_C;
    note_rom[46]   = HIGH_C;
    note_rom[47]   = HIGH_C;
    note_rom[48]   = MID_A;
    note_rom[49]   = MID_A;
    note_rom[50]   = MID_A;
    note_rom[51]   = MID_G;
    note_rom[52]   = MID_F;
    note_rom[53]   = MID_F;
    note_rom[54]   = MID_A;
    note_rom[55]   = MID_A;
    note_rom[56]   = MID_G;
    note_rom[57]   = MID_G;
    note_rom[58]   = MID_G;
    note_rom[59]   = MID_G;
    note_rom[60]   = MID_G;
    note_rom[61]   = MID_G;
    note_rom[62]   = SIL;;
    note_rom[63]   = MID_G;
    note_rom[64]   = MID_G;
    note_rom[65]   = MID_G;
    note_rom[66]   = MID_G;
    note_rom[67]   = MID_G;
    note_rom[68]   = MID_G;
    note_rom[69]   = MID_G;
    note_rom[70]   = MID_G;
    note_rom[71]   = MID_G;
    note_rom[72]   = MID_G;
    note_rom[73]   = MID_A;
    note_rom[74]   = MID_A;
    note_rom[75]   = MID_A;
    note_rom[76]   = MID_A;
    note_rom[77]   = MID_A;
    note_rom[78]   = MID_A;
    note_rom[79]   = MID_A;
    note_rom[80]   = MID_A;
    note_rom[81]   = MID_D;
    note_rom[82]   = MID_D;
    note_rom[83]   = MID_D;
    note_rom[84]   = MID_D;
    note_rom[85]   = MID_D;
    note_rom[86]   = MID_D;
    note_rom[87]   = MID_G;
    note_rom[88]   = MID_G;
    note_rom[89]   = MID_G;
    note_rom[90]   = MID_G;
    note_rom[91]   = MID_G;
    note_rom[92]   = MID_G;
    note_rom[93]   = MID_F;
    note_rom[94]   = MID_F;
    note_rom[95]   = MID_E;
    note_rom[96]   = MID_E;
    note_rom[97]   = MID_E;
    note_rom[98]   = MID_E;
    note_rom[99]   = LOW_G;
    note_rom[100]  = LOW_G;
    note_rom[101]  = LOW_G;
    note_rom[102]  = LOW_G;
    note_rom[103]  = MID_G;
    note_rom[104]  = MID_G;
    note_rom[105]  = MID_G;
    note_rom[106]  = MID_G;
    note_rom[107]  = MID_G;
    note_rom[108]  = MID_G;
    note_rom[109]  = MID_A;
    note_rom[110]  = MID_A;
    note_rom[111]  = MID_G;
    note_rom[112]  = MID_G;
    note_rom[113]  = MID_F;
    note_rom[114]  = MID_F;
    note_rom[115]  = MID_E;
    note_rom[116]  = MID_E;
    note_rom[117]  = MID_D;
    note_rom[118]  = MID_D;
    note_rom[119]  = MID_C;
    note_rom[120]  = MID_C;
    note_rom[121]  = MID_C;
    note_rom[122]  = MID_C;
    note_rom[123]  = MID_C;
    note_rom[124]  = MID_C;
    note_rom[125]  = MID_C;
    note_rom[126]  = MID_C;
    note_rom[127]  = MID_C;
    note_rom[128]  = MID_C;
    note_rom[129]  = MID_C;
    note_rom[130]  = LOW_G;
    note_rom[131]  = MID_E;
    note_rom[132]  = MID_E;
    note_rom[133]  = MID_E;
    note_rom[134]  = MID_E;
    note_rom[135]  = MID_E;
    note_rom[136]  = MID_E;
    note_rom[137]  = MID_E;
    note_rom[138]  = MID_E;
    note_rom[139]  = MID_E;
    note_rom[140]  = MID_E;
    note_rom[141]  = SIL;
    note_rom[142]  = MID_E;
    note_rom[143]  = MID_E;
    note_rom[144]  = MID_E;
    note_rom[145]  = MID_C;
    note_rom[146]  = MID_A;
    note_rom[147]  = MID_A;
    note_rom[148]  = MID_A;
    note_rom[149]  = MID_A;
    note_rom[150]  = MID_A;
    note_rom[151]  = MID_A;
    note_rom[152]  = MID_A;
    note_rom[153]  = MID_A;
    note_rom[154]  = MID_A;
    note_rom[155]  = SIL;
    note_rom[156]  = LOW_A;
    note_rom[157]  = LOW_A;
    note_rom[158]  = LOW_A;
    note_rom[159]  = LOW_A;
    note_rom[160]  = LOW_A;
    note_rom[161]  = LOW_A;
    note_rom[162]  = LOW_A;
    note_rom[163]  = LOW_A;
    note_rom[164]  = MID_D;
    note_rom[165]  = MID_D;
    note_rom[166]  = MID_D;
    note_rom[167]  = MID_D;
    note_rom[168]  = MID_D;
    note_rom[169]  = MID_D;
    note_rom[170]  = MID_E;
    note_rom[171]  = MID_D;
    note_rom[172]  = MID_D;
    note_rom[173]  = MID_C;
    note_rom[174]  = MID_C;
    note_rom[175]  = LOW_B;
    note_rom[176]  = LOW_B;
    note_rom[177]  = LOW_A;
    note_rom[178]  = LOW_A;
    note_rom[179]  = LOW_G;
    note_rom[180]  = LOW_G;
    note_rom[181]  = LOW_G;
    note_rom[182]  = LOW_G;
    note_rom[183]  = LOW_G;
    note_rom[184]  = LOW_G;
    note_rom[185]  = LOW_G;
    note_rom[186]  = LOW_G;
    note_rom[187]  = MID_C;
    note_rom[188]  = MID_C;
    note_rom[189]  = MID_C;
    note_rom[190]  = MID_C;
    note_rom[191]  = LOW_G;
    note_rom[192]  = LOW_G;
    note_rom[193]  = LOW_G;
    note_rom[194]  = LOW_G;
    note_rom[195]  = LOW_A;
    note_rom[196]  = LOW_A;
    note_rom[197]  = LOW_A;
    note_rom[198]  = LOW_A;
    note_rom[199]  = LOW_A;
    note_rom[200]  = LOW_A;
    note_rom[201]  = LOW_G;
    note_rom[202]  = LOW_G;
    note_rom[203]  = MID_C;
    note_rom[204]  = MID_C;
    note_rom[205]  = MID_C;
    note_rom[206]  = MID_C;
    note_rom[207]  = MID_D;
    note_rom[208]  = MID_D;
    note_rom[209]  = MID_D;
    note_rom[210]  = MID_D;
    note_rom[211]  = MID_E;
    note_rom[212]  = MID_E;
    note_rom[213]  = MID_E;
    note_rom[214]  = MID_E;
    note_rom[215]  = MID_E;
    note_rom[216]  = SIL;
    note_rom[217]  = MID_D;
    note_rom[218]  = MID_D;
    note_rom[219]  = MID_D;
    note_rom[220]  = MID_D;
    note_rom[221]  = MID_D;
    note_rom[222]  = MID_A;
    note_rom[223]  = MID_A;
    note_rom[224]  = MID_A;
    note_rom[225]  = MID_A;
    note_rom[226]  = MID_G;
    note_rom[227]  = MID_G;
    note_rom[228]  = MID_G;
    note_rom[229]  = MID_G;
    note_rom[230]  = MID_G;
    note_rom[231]  = MID_G;
    note_rom[232]  = MID_E;
    note_rom[233]  = MID_E;
    note_rom[234]  = MID_D;
    note_rom[235]  = MID_D;
    note_rom[236]  = MID_D;
    note_rom[237]  = MID_D;
    note_rom[238]  = MID_A;
    note_rom[239]  = MID_A;
    note_rom[240]  = MID_A;
    note_rom[241]  = MID_A;
    note_rom[242]  = MID_G;
    note_rom[243]  = MID_G;
    note_rom[244]  = MID_G;
    note_rom[245]  = MID_G;
    note_rom[246]  = SIL;
    note_rom[247]  = HIGH_C;
    note_rom[248]  = HIGH_C;
    note_rom[249]  = HIGH_C;
    note_rom[250]  = HIGH_C;
    note_rom[251]  = HIGH_C;
    note_rom[252]  = SIL;
    note_rom[253]  = HIGH_C;
    note_rom[254]  = HIGH_C;
    note_rom[255]  = MID_G;
    note_rom[256]  = MID_G;
    note_rom[257]  = MID_A;
    note_rom[258]  = MID_A;
    note_rom[259]  = MID_A;
    note_rom[260]  = MID_A;
    note_rom[261]  = MID_A;
    note_rom[262]  = MID_A;
    note_rom[263]  = HIGH_C;
    note_rom[264]  = HIGH_C;
    note_rom[265]  = MID_A;
    note_rom[266]  = MID_A;
    note_rom[267]  = MID_A;
    note_rom[268]  = MID_G;
    note_rom[269]  = MID_F;
    note_rom[270]  = MID_F;
    note_rom[271]  = MID_A;
    note_rom[272]  = MID_A;
    note_rom[273]  = MID_G;
    note_rom[274]  = MID_G;
    note_rom[275]  = MID_G;
    note_rom[276]  = MID_G;
    note_rom[277]  = MID_G;
    note_rom[278]  = SIL;
    note_rom[279]  = LOW_C;
    note_rom[280]  = LOW_C;
    note_rom[281]  = LOW_C;
    note_rom[282]  = LOW_C;
    note_rom[283]  = SIL;
    note_rom[284]  = LOW_C;
    note_rom[285]  = LOW_C;
    note_rom[286]  = LOW_C;
    note_rom[287]  = LOW_C;
    note_rom[288]  = MID_G;
    note_rom[289]  = MID_G;
    note_rom[290]  = MID_G;
    note_rom[291]  = MID_G;
    note_rom[292]  = MID_G;
    note_rom[293]  = MID_G;
    note_rom[294]  = MID_A;
    note_rom[295]  = MID_A;
    note_rom[296]  = MID_G;
    note_rom[297]  = MID_G;
    note_rom[298]  = MID_F;
    note_rom[299]  = MID_F;
    note_rom[300]  = MID_E;
    note_rom[301]  = MID_E;
    note_rom[302]  = MID_D;
    note_rom[303]  = MID_D;
    note_rom[304]  = MID_C;
    note_rom[305]  = MID_C;
    note_rom[306]  = MID_C;
    note_rom[307]  = MID_C;
    note_rom[308]  = LOW_G;
    note_rom[309]  = LOW_G;
    note_rom[310]  = LOW_G;
    note_rom[311]  = LOW_G;
    note_rom[312]  = MID_C;
    note_rom[313]  = MID_C;
    note_rom[314]  = MID_C;
    note_rom[315]  = MID_C;
    note_rom[316]  = LOW_G;
    note_rom[317]  = LOW_G;
    note_rom[318]  = LOW_G;
    note_rom[319]  = LOW_G;
    note_rom[320]  = MID_E;
    note_rom[321]  = MID_E;
    note_rom[322]  = MID_E;
    note_rom[323]  = MID_E;
    note_rom[324]  = MID_C;
    note_rom[325]  = MID_C;
    note_rom[326]  = MID_C;
    note_rom[327]  = MID_C;
    note_rom[328]  = MID_G;
    note_rom[329]  = MID_G;
    note_rom[330]  = MID_G;
    note_rom[331]  = MID_G;
    note_rom[332]  = MID_G;
    note_rom[333]  = MID_A;
    note_rom[334]  = MID_A;
    note_rom[335]  = MID_A;
    note_rom[336]  = MID_G;
    note_rom[337]  = MID_G;
    note_rom[338]  = MID_G;
    note_rom[339]  = MID_G;
    note_rom[340]  = SIL;
    note_rom[341]  = MID_G;
    note_rom[342]  = MID_G;
    note_rom[343]  = MID_G;
    note_rom[344]  = MID_G;
    note_rom[345]  = MID_G;
    note_rom[346]  = MID_G;
    note_rom[347]  = HIGH_C;
    note_rom[348]  = HIGH_C;
    note_rom[349]  = HIGH_C;
    note_rom[350]  = HIGH_C;
    note_rom[351]  = HIGH_C;
    note_rom[352]  = HIGH_C;
    note_rom[353]  = HIGH_C;
    note_rom[354]  = HIGH_C;
    note_rom[355]  = HIGH_C;
    note_rom[356]  = MID_A;
    note_rom[357]  = MID_A;
    note_rom[358]  = MID_A;
    note_rom[359]  = MID_G;
    note_rom[360]  = MID_F;
    note_rom[361]  = MID_F;
    note_rom[362]  = MID_A;
    note_rom[363]  = MID_A;
    note_rom[364]  = MID_G;
    note_rom[365]  = MID_G;
    note_rom[366]  = MID_G;
    note_rom[367]  = MID_G;
    note_rom[368]  = SIL;
    note_rom[369]  = MID_G;
    note_rom[370]  = MID_G;
    note_rom[371]  = MID_G;
    note_rom[372]  = MID_G;
    note_rom[373]  = MID_G;
    note_rom[374]  = MID_G;
    note_rom[375]  = MID_G;
    note_rom[376]  = MID_G;
    note_rom[377]  = MID_G;
    note_rom[378]  = MID_G;
    note_rom[379]  = MID_G;
    note_rom[380]  = MID_G;
    note_rom[381]  = MID_A;
    note_rom[382]  = MID_A;
    note_rom[383]  = MID_A;
    note_rom[384]  = MID_A;
    note_rom[385]  = MID_A;
    note_rom[386]  = MID_A;
    note_rom[387]  = MID_A;
    note_rom[388]  = MID_A;
    note_rom[389]  = MID_D;
    note_rom[390]  = MID_D;
    note_rom[391]  = MID_D;
    note_rom[392]  = MID_D;
    note_rom[393]  = MID_D;
    note_rom[394]  = MID_D;
    note_rom[395]  = MID_G;
    note_rom[396]  = MID_G;
    note_rom[397]  = MID_G;
    note_rom[398]  = MID_G;
    note_rom[399]  = MID_G;
    note_rom[400]  = MID_G;
    note_rom[401]  = MID_F;
    note_rom[402]  = MID_F;
    note_rom[403]  = MID_E;
    note_rom[404]  = MID_E;
    note_rom[405]  = MID_E;
    note_rom[406]  = MID_E;
    note_rom[407]  = LOW_G;
    note_rom[408]  = LOW_G;
    note_rom[409]  = LOW_G;
    note_rom[410]  = LOW_G;
    note_rom[411]  = MID_G;
    note_rom[412]  = MID_G;
    note_rom[413]  = MID_G;
    note_rom[414]  = MID_G;
    note_rom[415]  = MID_G;
    note_rom[416]  = MID_G;
    note_rom[417]  = MID_A;
    note_rom[418]  = MID_A;
    note_rom[419]  = MID_G;
    note_rom[420]  = MID_G;
    note_rom[421]  = MID_F;
    note_rom[422]  = MID_F;
    note_rom[423]  = MID_E;
    note_rom[424]  = MID_E;
    note_rom[425]  = MID_D;
    note_rom[426]  = MID_D;
    note_rom[427]  = MID_C;
    note_rom[428]  = MID_C;
    note_rom[429]  = MID_C;
    note_rom[430]  = MID_C;
    note_rom[431]  = MID_C;
    note_rom[432]  = MID_C;
    note_rom[433]  = MID_C;
    note_rom[434]  = MID_C;
    note_rom[435]  = MID_C;
    note_rom[436]  = MID_C;
    note_rom[437]  = MID_C;
    note_rom[438]  = LOW_G;
    note_rom[439]  = MID_E;
    note_rom[440]  = MID_E;
    note_rom[441]  = MID_E;
    note_rom[442]  = MID_E;
    note_rom[443]  = MID_E;
    note_rom[444]  = MID_E;
    note_rom[445]  = MID_E;
    note_rom[446]  = MID_E;
    note_rom[447]  = MID_E;
    note_rom[448]  = MID_E;
    note_rom[449]  = SIL;
    note_rom[450]  = MID_E;
    note_rom[451]  = MID_E;
    note_rom[452]  = MID_E;
    note_rom[453]  = MID_C;
    note_rom[454]  = MID_A;
    note_rom[455]  = MID_A;
    note_rom[456]  = MID_A;
    note_rom[457]  = MID_A;
    note_rom[458]  = MID_A;
    note_rom[459]  = MID_A;
    note_rom[460]  = MID_A;
    note_rom[461]  = MID_A;
    note_rom[462]  = MID_A;
    note_rom[463]  = SIL;
    note_rom[464]  = LOW_A;
    note_rom[465]  = LOW_A;
    note_rom[466]  = LOW_A;
    note_rom[467]  = LOW_A;
    note_rom[468]  = LOW_A;
    note_rom[469]  = LOW_A;
    note_rom[470]  = LOW_A;
    note_rom[471]  = LOW_A;
    note_rom[472]  = MID_D;
    note_rom[473]  = MID_D;
    note_rom[474]  = MID_D;
    note_rom[475]  = MID_D;
    note_rom[476]  = MID_D;
    note_rom[477]  = MID_D;
    note_rom[478]  = MID_E;
    note_rom[479]  = MID_D;
    note_rom[480]  = MID_D;
    note_rom[481]  = MID_C;
    note_rom[482]  = MID_C;
    note_rom[483]  = LOW_B;
    note_rom[484]  = LOW_B;
    note_rom[485]  = LOW_A;
    note_rom[486]  = LOW_A;
    note_rom[487]  = LOW_G;
    note_rom[488]  = LOW_G;
    note_rom[489]  = LOW_G;
    note_rom[490]  = LOW_G;
    note_rom[491]  = LOW_G;
    note_rom[492]  = LOW_G;
    note_rom[493]  = LOW_G;
    note_rom[494]  = LOW_G;
    note_rom[495]  = MID_C;
    note_rom[496]  = MID_C;
    note_rom[497]  = MID_C;
    note_rom[498]  = MID_C;
    note_rom[499]  = LOW_G;
    note_rom[500]  = LOW_G;
    note_rom[501]  = LOW_G;
    note_rom[502]  = LOW_G;
    note_rom[503]  = LOW_A;
    note_rom[504]  = LOW_A;
    note_rom[505]  = LOW_A;
    note_rom[506]  = LOW_A;
    note_rom[507]  = LOW_A;
    note_rom[508]  = LOW_A;
    note_rom[509]  = LOW_G;
    note_rom[510]  = LOW_G;
    note_rom[511]  = MID_C;


 //Call of Silence   
    // ====== 第二首歌(地址 512-1023) ======
    note_rom[512] = MID_D;
    note_rom[513] = MID_D;
    note_rom[514] = MID_A;
    note_rom[515] = MID_A;
    note_rom[516] = MID_A;
    note_rom[517] = MID_A;
    note_rom[518] = MID_A;
    note_rom[519] = MID_A;
    note_rom[520] = MID_A;
    note_rom[521] = MID_A;
    note_rom[522] = MID_A;
    note_rom[523] = MID_E;
    note_rom[524] = MID_E;
    note_rom[525] = MID_E;
    note_rom[526] = MID_E;
    note_rom[527] = MID_E;
    note_rom[528] = MID_E;
    note_rom[529] = MID_E;
    note_rom[530] = MID_D;
    note_rom[531] = MID_F;
    note_rom[532] = MID_F;
    note_rom[533] = MID_F;
    note_rom[534] = MID_F;
    note_rom[535] = MID_F;
    note_rom[536] = MID_F;
    note_rom[537] = MID_F;
    note_rom[538] = MID_F;
    note_rom[539] = MID_F;
    note_rom[540] = SIL;
    note_rom[541] = MID_D;
    note_rom[542] = MID_D;
    note_rom[543] = MID_A;
    note_rom[544] = MID_A;
    note_rom[545] = MID_A;
    note_rom[546] = MID_A;
    note_rom[547] = MID_A;
    note_rom[548] = MID_A;
    note_rom[549] = MID_A;
    note_rom[550] = MID_A;
    note_rom[551] = HIGH_E;
    note_rom[552] = HIGH_E;
    note_rom[553] = HIGH_E;
    note_rom[554] = HIGH_E;
    note_rom[555] = HIGH_E;
    note_rom[556] = HIGH_E;
    note_rom[557] = HIGH_E;
    note_rom[558] = HIGH_A;
    note_rom[559] = HIGH_A;
    note_rom[560] = HIGH_A;
    note_rom[561] = HIGH_A;
    note_rom[562] = HIGH_A;
    note_rom[563] = HIGH_A;
    note_rom[564] = HIGH_A;
    note_rom[565] = HIGH_A;
    note_rom[566] = HIGH_A;
    note_rom[567] = HIGH_A;
    note_rom[568] = HIGH_A;
    note_rom[569] = HIGH_A;
    note_rom[570] = HIGH_A;
    note_rom[571] = HIGH_E;
    note_rom[572] = HIGH_E;
    note_rom[573] = HIGH_E;
    note_rom[574] = HIGH_E;
    note_rom[575] = HIGH_E;
    note_rom[576] = HIGH_E;
    note_rom[577] = HIGH_E;
    note_rom[578] = HIGH_E;
    note_rom[579] = HIGH_F;
    note_rom[580] = HIGH_C;
    note_rom[581] = HIGH_C;
    note_rom[582] = HIGH_C;
    note_rom[583] = HIGH_C;
    note_rom[584] = HIGH_C;
    note_rom[585] = HIGH_C;
    note_rom[586] = HIGH_C;
    note_rom[587] = HIGH_C;
    note_rom[588] = HIGH_C;
    note_rom[589] = SIL;
    note_rom[590] = HIGH_C;
    note_rom[591] = HIGH_C;
    note_rom[592] = MID_A;
    note_rom[593] = HIGH_C;
    note_rom[594] = HIGH_C;
    note_rom[595] = HIGH_C;
    note_rom[596] = HIGH_C;
    note_rom[597] = HIGH_C;
    note_rom[598] = HIGH_C;
    note_rom[599] = HIGH_C;
    note_rom[600] = SIL;
    note_rom[601] = HIGH_G;
    note_rom[602] = HIGH_G;
    note_rom[603] = HIGH_F;
    note_rom[604] = HIGH_G;
    note_rom[605] = HIGH_G;
    note_rom[606] = HIGH_G;
    note_rom[607] = HIGH_G;
    note_rom[608] = HIGH_G;
    note_rom[609] = HIGH_G;
    note_rom[610] = HIGH_G;
    note_rom[611] = HIGH_F;
    note_rom[612] = HIGH_D;
    note_rom[613] = HIGH_D;
    note_rom[614] = HIGH_D;
    note_rom[615] = HIGH_D;
    note_rom[616] = HIGH_D;
    note_rom[617] = SIL;
    note_rom[618] = SIL;
    note_rom[619] = HIGH_A;
    note_rom[620] = HIGH_A;
    note_rom[621] = HIGH_G;
    note_rom[622] = HIGH_G;
    note_rom[623] = HIGH_G;
    note_rom[624] = HIGH_G;
    note_rom[625] = HIGH_F;
    note_rom[626] = HIGH_F;
    note_rom[627] = HIGH_F;
    note_rom[628] = HIGH_F;
    note_rom[629] = HIGH_C;
    note_rom[630] = HIGH_C;
    note_rom[631] = HIGH_F;
    note_rom[632] = HIGH_F;
    note_rom[633] = HIGH_F;
    note_rom[634] = HIGH_F;
    note_rom[635] = HIGH_E;
    note_rom[636] = HIGH_E;
    note_rom[637] = HIGH_F;
    note_rom[638] = HIGH_F;
    note_rom[639] = HIGH_F;
    note_rom[640] = HIGH_F;
    note_rom[641] = SIL;
    note_rom[642] = HIGH_A;
    note_rom[643] = HIGH_A;
    note_rom[644] = HIGH_G;
    note_rom[645] = HIGH_G;
    note_rom[646] = HIGH_G;
    note_rom[647] = HIGH_G;
    note_rom[648] = HIGH_F;
    note_rom[649] = HIGH_F;
    note_rom[650] = HIGH_F;
    note_rom[651] = HIGH_F;
    note_rom[652] = HIGH_A;
    note_rom[653] = HIGH_A;
    note_rom[654] = HIGH_F;
    note_rom[655] = HIGH_F;
    note_rom[656] = HIGH_F;
    note_rom[657] = HIGH_F;
    note_rom[658] = SIL;
    note_rom[659] = HIGH_F;
    note_rom[660] = HIGH_F;
    note_rom[661] = HIGH_E;
    note_rom[662] = HIGH_E;
    note_rom[663] = MID_A;
    note_rom[664] = HIGH_D;
    note_rom[665] = HIGH_D;
    note_rom[666] = HIGH_D;
    note_rom[667] = HIGH_D;
    note_rom[668] = HIGH_D;
    note_rom[669] = HIGH_D;
    note_rom[670] = HIGH_D;
    note_rom[671] = HIGH_D;
    note_rom[672] = HIGH_E;
    note_rom[673] = HIGH_E;
    note_rom[674] = HIGH_E;
    note_rom[675] = HIGH_E;
    note_rom[676] = HIGH_E;
    note_rom[677] = HIGH_E;
    note_rom[678] = HIGH_E;
    note_rom[679] = HIGH_G;
    note_rom[680] = HIGH_F;
    note_rom[681] = HIGH_F;
    note_rom[682] = HIGH_F;
    note_rom[683] = HIGH_F;
    note_rom[684] = HIGH_F;
    note_rom[685] = HIGH_F;
    note_rom[686] = HIGH_F;
    note_rom[687] = HIGH_F;
    note_rom[688] = HIGH_F;
    note_rom[689] = SIL;
    note_rom[690] = HIGH_F;
    note_rom[691] = HIGH_F;
    note_rom[692] = HIGH_E;
    note_rom[693] = HIGH_E;
    note_rom[694] = MID_A;
    note_rom[695] = HIGH_D;
    note_rom[696] = HIGH_D;
    note_rom[697] = HIGH_D;
    note_rom[698] = HIGH_D;
    note_rom[699] = HIGH_D;
    note_rom[700] = HIGH_D;
    note_rom[701] = SIL;
    note_rom[702] = SIL;
    note_rom[703] = HIGH_A;
    note_rom[704] = HIGH_A;
    note_rom[705] = HIGH_G;
    note_rom[706] = HIGH_G;
    note_rom[707] = HIGH_G;
    note_rom[708] = HIGH_G;
    note_rom[709] = HIGH_F;
    note_rom[710] = HIGH_F;
    note_rom[711] = HIGH_F;
    note_rom[712] = HIGH_F;
    note_rom[713] = HIGH_C2;
    note_rom[714] = HIGH_C2;
    note_rom[715] = HIGH_C2;
    note_rom[716] = HIGH_C2;
    note_rom[717] = HIGH_C2;
    note_rom[718] = HIGH_C2;
    note_rom[719] = HIGH_G;
    note_rom[720] = HIGH_G;
    note_rom[721] = HIGH_F;
    note_rom[722] = HIGH_F;
    note_rom[723] = HIGH_F;
    note_rom[724] = HIGH_F;
    note_rom[725] = HIGH_F;
    note_rom[726] = HIGH_F;
    note_rom[727] = SIL;
    note_rom[728] = HIGH_D;
    note_rom[729] = HIGH_D;
    note_rom[730] = HIGH_F;
    note_rom[731] = HIGH_F;
    note_rom[732] = HIGH_G;
    note_rom[733] = HIGH_G;
    note_rom[734] = HIGH_G;
    note_rom[735] = HIGH_G;
    note_rom[736] = HIGH_G;
    note_rom[737] = HIGH_G;
    note_rom[738] = HIGH_F;
    note_rom[739] = HIGH_F;
    note_rom[740] = HIGH_G;
    note_rom[741] = HIGH_G;
    note_rom[742] = HIGH_A;
    note_rom[743] = HIGH_A;
    note_rom[744] = HIGH_G;
    note_rom[745] = HIGH_G;
    note_rom[746] = HIGH_G;
    note_rom[747] = HIGH_G;
    note_rom[748] = HIGH_G;
    note_rom[749] = HIGH_F;
    note_rom[750] = HIGH_F;
    note_rom[751] = HIGH_F;
    note_rom[752] = HIGH_F;
    note_rom[753] = HIGH_F;
    note_rom[754] = HIGH_F;
    note_rom[755] = SIL;
    note_rom[756] = HIGH_F;
    note_rom[757] = HIGH_F;
    note_rom[758] = HIGH_E;
    note_rom[759] = HIGH_E;
    note_rom[760] = MID_A;
    note_rom[761] = HIGH_D;
    note_rom[762] = HIGH_D;
    note_rom[763] = HIGH_D;
    note_rom[764] = HIGH_D;
    note_rom[765] = HIGH_D;
    note_rom[766] = HIGH_D;
    note_rom[767] = HIGH_D;
    note_rom[768] = HIGH_D;
    note_rom[769] = HIGH_E;
    note_rom[770] = HIGH_E;
    note_rom[771] = HIGH_E;
    note_rom[772] = HIGH_E;
    note_rom[773] = HIGH_E;
    note_rom[774] = HIGH_E;
    note_rom[775] = HIGH_E;
    note_rom[776] = HIGH_G;
    note_rom[777] = HIGH_F;
    note_rom[778] = HIGH_F;
    note_rom[779] = HIGH_F;
    note_rom[780] = HIGH_F;
    note_rom[781] = HIGH_F;
    note_rom[782] = HIGH_F;
    note_rom[783] = HIGH_F;
    note_rom[784] = HIGH_F;
    note_rom[785] = HIGH_F;
    note_rom[786] = SIL;
    note_rom[787] = HIGH_F;
    note_rom[788] = HIGH_F;
    note_rom[789] = HIGH_E;
    note_rom[790] = HIGH_E;
    note_rom[791] = MID_A;
    note_rom[792] = HIGH_D;
    note_rom[793] = HIGH_D;
    note_rom[794] = HIGH_D;
    note_rom[795] = HIGH_D;
    note_rom[796] = HIGH_D;
    note_rom[797] = HIGH_D;
    note_rom[798] = SIL;
    note_rom[799] = SIL;
    note_rom[800] = HIGH_A;
    note_rom[801] = HIGH_A;
    note_rom[802] = HIGH_G;
    note_rom[803] = HIGH_G;
    note_rom[804] = HIGH_G;
    note_rom[805] = HIGH_G;
    note_rom[806] = HIGH_F;
    note_rom[807] = HIGH_F;
    note_rom[808] = HIGH_F;
    note_rom[809] = HIGH_F;
    note_rom[810] = HIGH_C2;
    note_rom[811] = HIGH_C2;
    note_rom[812] = HIGH_C2;
    note_rom[813] = HIGH_C2;
    note_rom[814] = HIGH_C2;
    note_rom[815] = HIGH_C2;
    note_rom[816] = HIGH_G;
    note_rom[817] = HIGH_G;
    note_rom[818] = HIGH_F;
    note_rom[819] = HIGH_F;
    note_rom[820] = HIGH_F;
    note_rom[821] = HIGH_F;
    note_rom[822] = HIGH_F;
    note_rom[823] = HIGH_F;
    note_rom[824] = SIL;
    note_rom[825] = HIGH_D;
    note_rom[826] = HIGH_D;
    note_rom[827] = HIGH_F;
    note_rom[828] = HIGH_F;
    note_rom[829] = HIGH_G;
    note_rom[830] = HIGH_G;
    note_rom[831] = HIGH_G;
    note_rom[832] = HIGH_G;
    note_rom[833] = HIGH_G;
    note_rom[834] = HIGH_G;
    note_rom[835] = HIGH_G;
    note_rom[836] = HIGH_F;
    note_rom[837] = HIGH_F;
    note_rom[838] = HIGH_G;
    note_rom[839] = HIGH_G;
    note_rom[840] = HIGH_A;
    note_rom[841] = HIGH_A;
    note_rom[842] = HIGH_G;
    note_rom[843] = HIGH_G;
    note_rom[844] = HIGH_G;
    note_rom[845] = HIGH_G;
    note_rom[846] = HIGH_G;
    note_rom[847] = HIGH_F;
    note_rom[848] = HIGH_F;
    note_rom[849] = HIGH_F;
    note_rom[850] = HIGH_F;
    note_rom[851] = HIGH_F;
    note_rom[852] = HIGH_F;
    note_rom[853] = SIL;
    note_rom[854] = HIGH_F;
    note_rom[855] = HIGH_F;
    note_rom[856] = HIGH_E;
    note_rom[857] = HIGH_E;
    note_rom[858] = MID_A;
    note_rom[859] = HIGH_D;
    note_rom[860] = HIGH_D;
    note_rom[861] = HIGH_D;
    note_rom[862] = HIGH_D;
    note_rom[863] = HIGH_D;
    note_rom[864] = HIGH_D;
    note_rom[865] = HIGH_D;
    note_rom[866] = HIGH_D;
    note_rom[867] = HIGH_E;
    note_rom[868] = HIGH_E;
    note_rom[869] = HIGH_E;
    note_rom[870] = HIGH_E;
    note_rom[871] = HIGH_E;
    note_rom[872] = HIGH_E;
    note_rom[873] = HIGH_E;
    note_rom[874] = HIGH_G;
    note_rom[875] = HIGH_F;
    note_rom[876] = HIGH_F;
    note_rom[877] = HIGH_F;
    note_rom[878] = HIGH_F;
    note_rom[879] = HIGH_F;
    note_rom[880] = HIGH_F;
    note_rom[881] = HIGH_F;
    note_rom[882] = HIGH_F;
    note_rom[883] = HIGH_F;
    note_rom[884] = SIL;
    note_rom[885] = HIGH_F;
    note_rom[886] = HIGH_F;
    note_rom[887] = HIGH_E;
    note_rom[888] = HIGH_E;
    note_rom[889] = MID_A;
    note_rom[890] = HIGH_D;
    note_rom[891] = HIGH_D;
    note_rom[892] = HIGH_D;
    note_rom[893] = HIGH_D;
    note_rom[894] = HIGH_D;
    note_rom[895] = HIGH_D;
    note_rom[896] = SIL;
    note_rom[897] = SIL;
    note_rom[898] = HIGH_A;
    note_rom[899] = HIGH_A;
    note_rom[900] = HIGH_G;
    note_rom[901] = HIGH_G;
    note_rom[902] = HIGH_G;
    note_rom[903] = HIGH_G;
    note_rom[904] = HIGH_F;
    note_rom[905] = HIGH_F;
    note_rom[906] = HIGH_F;
    note_rom[907] = HIGH_F;
    note_rom[908] = HIGH_C2;
    note_rom[909] = HIGH_C2;
    note_rom[910] = HIGH_C2;
    note_rom[911] = HIGH_C2;
    note_rom[912] = HIGH_C2;
    note_rom[913] = HIGH_C2;
    note_rom[914] = HIGH_G;
    note_rom[915] = HIGH_G;
    note_rom[916] = HIGH_F;
    note_rom[917] = HIGH_F;
    note_rom[918] = HIGH_F;
    note_rom[919] = HIGH_F;
    note_rom[920] = HIGH_F;
    note_rom[921] = HIGH_F;
    note_rom[922] = SIL;
    note_rom[923] = HIGH_D;
    note_rom[924] = HIGH_D;
    note_rom[925] = HIGH_F;
    note_rom[926] = HIGH_F;
    note_rom[927] = HIGH_G;
    note_rom[928] = HIGH_G;
    note_rom[929] = HIGH_G;
    note_rom[930] = HIGH_G;
    note_rom[931] = HIGH_G;
    note_rom[932] = HIGH_G;
    note_rom[933] = HIGH_G;
    note_rom[934] = HIGH_F;
    note_rom[935] = HIGH_F;
    note_rom[936] = HIGH_G;
    note_rom[937] = HIGH_G;
    note_rom[938] = HIGH_A;
    note_rom[939] = HIGH_A;
    note_rom[940] = HIGH_G;
    note_rom[941] = HIGH_G;
    note_rom[942] = HIGH_G;
    note_rom[943] = HIGH_G;
    note_rom[944] = HIGH_G;
    note_rom[945] = HIGH_F;
    note_rom[946] = HIGH_F;
    note_rom[947] = HIGH_F;
    note_rom[948] = HIGH_F;
    note_rom[949] = HIGH_F;
    note_rom[950] = HIGH_F;
    note_rom[951] = SIL;
    note_rom[952] = HIGH_F;
    note_rom[953] = HIGH_F;
    note_rom[954] = HIGH_E;
    note_rom[955] = HIGH_E;
    note_rom[956] = MID_A;
    note_rom[957] = HIGH_D;
    note_rom[958] = HIGH_D;
    note_rom[959] = HIGH_D;
    note_rom[960] = HIGH_D;
    note_rom[961] = HIGH_D;
    note_rom[962] = HIGH_D;
    note_rom[963] = HIGH_D;
    note_rom[964] = HIGH_D;
    note_rom[965] = HIGH_E;
    note_rom[966] = HIGH_E;
    note_rom[967] = HIGH_E;
    note_rom[968] = HIGH_E;
    note_rom[969] = HIGH_E;
    note_rom[970] = HIGH_E;
    note_rom[971] = HIGH_E;
    note_rom[972] = HIGH_G;
    note_rom[973] = HIGH_F;
    note_rom[974] = HIGH_F;
    note_rom[975] = HIGH_F;
    note_rom[976] = HIGH_F;
    note_rom[977] = HIGH_F;
    note_rom[978] = HIGH_F;
    note_rom[979] = HIGH_F;
    note_rom[980] = HIGH_F;
    note_rom[981] = HIGH_F;
    note_rom[982] = SIL;
    note_rom[983] = HIGH_F;
    note_rom[984] = HIGH_F;
    note_rom[985] = HIGH_E;
    note_rom[986] = HIGH_E;
    note_rom[987] = MID_A;
    note_rom[988] = HIGH_D;
    note_rom[989] = HIGH_D;
    note_rom[990] = HIGH_D;
    note_rom[991] = HIGH_D;
    note_rom[992] = HIGH_D;
    note_rom[993] = HIGH_D;
    note_rom[994] = SIL;
    note_rom[995] = SIL;
    note_rom[996] = HIGH_A;
    note_rom[997] = HIGH_A;
    note_rom[998] = HIGH_G;
    note_rom[999] = HIGH_G;
    note_rom[1000] = HIGH_G;
    note_rom[1001] = HIGH_G;
    note_rom[1002] = HIGH_F;
    note_rom[1003] = HIGH_F;
    note_rom[1004] = HIGH_F;
    note_rom[1005] = HIGH_F;
    note_rom[1006] = HIGH_C2;
    note_rom[1007] = HIGH_C2;
    note_rom[1008] = HIGH_C2;
    note_rom[1009] = HIGH_C2;
    note_rom[1010] = HIGH_C2;
    note_rom[1011] = HIGH_C2;
    note_rom[1012] = HIGH_G;
    note_rom[1013] = HIGH_G;
    note_rom[1014] = HIGH_F;
    note_rom[1015] = HIGH_F;
    note_rom[1016] = HIGH_F;
    note_rom[1017] = HIGH_F;
    note_rom[1018] = HIGH_F;
    note_rom[1019] = HIGH_F;
    note_rom[1020] = SIL;
    note_rom[1021] = HIGH_D;
    note_rom[1022] = HIGH_D;
    note_rom[1023] = HIGH_F;

    // ... 添加更多音 MID_A;符直到地址1023 ...
  end

  always @ (posedge clk, negedge rst_n) begin
    if (rst_n == 1'b0)
      music <= SIL;
    else
      music <= note_rom[cnt]; // 直接ROM查找
  end

endmodule